module test (
     output   [5:0]out
	      );
			
	wire   [5:0]a;
	assign a = 3;
	assign out = a;
	
	
endmodule
	